`define DELAY 10
module alu32_tb();

wire [31:0] R;
wire Zero,Overflow;
reg [31:0] A;
reg [31:0] B;
reg [2:0] Op; 


alu32 u1( R, A, B, Op, Zero,Overflow);

initial begin

// AND Tests
A = 32'b11100001100000001101001110000101;
B = 32'b11100000000111000000001110000010;
Op = 3'b000;
#`DELAY;
A = 32'b11010101101011001011010100101010;
B = 32'b01011110001100000001110011110110;
Op = 3'b000;
#`DELAY;
A = 32'b10101010101010101010101010101010;
B = 32'b01010101010101010101010101010101;
Op = 3'b000;
#`DELAY;


//OR Tests
A = 32'b11100000000000001111111111111111;
B = 32'b00000011100000001111111000001111;
Op = 3'b001;
#`DELAY;
A = 32'b11010101101011001011010100101010;
B = 32'b01011110001100000001110011110110;
Op = 3'b001;
#`DELAY;
A = 32'b10101010101010101010101010101010;
B = 32'b01010101010101010101010101010101;
Op = 3'b001;
#`DELAY;

//ADD Tests
// Overflow 
A = 32'b01000000000000000000000000000000; 
B = 32'b01000000000000000000000000000000;
Op = 3'b010;
#`DELAY;
// 12 + 17 = 29
A = 32'b00000000000000000000000000001100; 
B = 32'b00000000000000000000000000010001;
Op = 3'b010;
#`DELAY;
// 174 + 13 = 187
A = 32'b00000000000000000000000010101110; 
B = 32'b00000000000000000000000000001101;
Op = 3'b010;
#`DELAY;


//XOR Tests
A = 32'b11100000000000001111111111111111;
B = 32'b00000011100000001111111000001111;
Op = 3'b011;
#`DELAY;
A = 32'b11010101101011001011010100101010;
B = 32'b01011110001100000001110011110110;
Op = 3'b011;
#`DELAY;
A = 32'b10101010101010101010101010101010;
B = 32'b01010101010101010101010101010101;
Op = 3'b011;
#`DELAY;


//SUB Tests
// Overflow
A = 32'b00000000000000000000000000100000; 
B = 32'b10000000000000000000000000011001;
Op = 3'b100;
#`DELAY;
// 17 - 12 = 5
A = 32'b00000000000000000000000000010001;
B = 32'b00000000000000000000000000001100;
Op = 3'b100;
#`DELAY;
// 174 - 13 = 161
A = 32'b00000000000000000000000010101110; 
B = 32'b00000000000000000000000000001101;
Op = 3'b100;
#`DELAY;

//Arithmetic Right Shift
A = 32'b11111000000000000000000000011111;
B = 32'b00000000000000000000000000000101;
Op = 3'b101;
#`DELAY;
A = 32'b00011100011100000000001111000111;
B = 32'b00000000000000000000000000000111;
Op = 3'b101;
#`DELAY;
A = 32'b10101010101010101010101010101010;
B = 32'b00000000000000000000000000011111;
Op = 3'b101;
#`DELAY;


// Logic Left Shift
A = 32'b11111000000000000000000000010011;
B = 32'b00000000000000000000000000000101;
Op = 3'b110;
#`DELAY;
A = 32'b00011100011100000000001111000111;
B = 32'b00000000000000000000000000000111;
Op = 3'b110;
#`DELAY;
A = 32'b01010100101010101010101010101010;
B = 32'b00000000000000000000000000011111;
Op = 3'b110;
#`DELAY;

//NOR Tests
A = 32'b11100000000000001111111111111111;
B = 32'b00000011100000001111111000001111;
Op = 3'b111;
#`DELAY;
A = 32'b11010101101011001011010100101010;
B = 32'b01011110001100000001110011110110;
Op = 3'b111;
#`DELAY;
A = 32'b10101010101010101010101010101010;
B = 32'b01010101010101010101010101010101;
Op = 3'b111;

end

initial
begin
$monitor("time = %2d, A = %32b, B = %32b, Operation = %3b, Result = %32b, Zero=%1b, Overflow=%1b", $time, A, B, Op, R, Zero,Overflow);
end

endmodule